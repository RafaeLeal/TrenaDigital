library IEEE;
use IEEE.Std_logic_1164.all;
use IEEE.Std_logic_arith.all;
use ieee.std_logic_unsigned.all;
ENTITY SD_sensor_de_distancia IS
PORT (
		CLK 			: IN STD_LOGIC;
		CLK2 			: IN STD_LOGIC;
		LIGA 			: IN STD_LOGIC;
		MEDIR 			: IN STD_LOGIC;
		ECHO 			: IN STD_LOGIC;
		RESET 			: IN STD_LOGIC;
		MEDIDA 			: OUT STD_LOGIC_VECTOR(15 downto 0);
		PRONTO 			: OUT STD_LOGIC;
		TRIGGER 		: OUT STD_LOGIC;
		UC_DEBUG_ESTADO : OUT STD_LOGIC_VECTOR(2 downto 0);
		A7SEG3 			: OUT STD_LOGIC_VECTOR(6 downto 0);
		A7SEG2 			: OUT STD_LOGIC_VECTOR(6 downto 0);
		A7SEG1 			: OUT STD_LOGIC_VECTOR(6 downto 0);
		A7SEG0 			: OUT STD_LOGIC_VECTOR(6 downto 0);
		SERIAL 			: OUT STD_LOGIC;
		MODO_ATUAL 		: OUT STD_LOGIC;
		CLK2_OUT 		: OUT STD_LOGIC
);
END ENTITY;
ARCHITECTURE arch_SD_sensor_de_distancia OF SD_sensor_de_distancia IS

COMPONENT UC_sensor_de_distancia
PORT(
	CLK : IN STD_LOGIC;
	MEDIR : IN STD_LOGIC;
	ECHO : IN STD_LOGIC;
	RESET : IN STD_LOGIC;
	TRIGGER : OUT STD_LOGIC;
	PRONTO : OUT STD_LOGIC;
	DEBUG_ESTADO : OUT STD_LOGIC_VECTOR(2 downto 0)
);
END COMPONENT;
COMPONENT FD_sensor_de_distancia
PORT(
	CLK : IN STD_LOGIC;
	ECHO : IN STD_LOGIC;
	RESET : IN STD_LOGIC;
	MEDIDA : OUT STD_LOGIC_VECTOR(15 downto 0);
	A7SEG3 : OUT STD_LOGIC_VECTOR(6 downto 0);
	A7SEG2 : OUT STD_LOGIC_VECTOR(6 downto 0);
	A7SEG1 : OUT STD_LOGIC_VECTOR(6 downto 0);
	A7SEG0 : OUT STD_LOGIC_VECTOR(6 downto 0);
	SAIDA_SERIAL : OUT STD_LOGIC
	);
END COMPONENT;
SIGNAL MEDIR_LIGADO : STD_LOGIC;

BEGIN
MEDIR_LIGADO <= MEDIR AND LIGA;
MODO_ATUAL <= LIGA;
CLK2_OUT <= CLK;
FLUXO_DE_DADOS: FD_sensor_de_distancia PORT MAP (
	CLK,
	ECHO,
	RESET,
	MEDIDA,
	A7SEG3,
	A7SEG2,
	A7SEG1,
	A7SEG0,
	SERIAL
	);
UNIDADE_DE_CONTROLE : UC_sensor_de_distancia PORT MAP (
	CLK,
	MEDIR_LIGADO,
	ECHO,
	RESET,
	TRIGGER,
	PRONTO,
	UC_DEBUG_ESTADO
	);
	
-- TODO PORT MAPPING
END ARCHITECTURE;